
module clock50to25 (
	clk_in_clk,
	reset_reset,
	clk_out_clk);	

	input		clk_in_clk;
	input		reset_reset;
	output		clk_out_clk;
endmodule
