-- clock50to150.vhd

-- Generated using ACDS version 23.1 991

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity clock50to150 is
	port (
		clk_in_clk  : in  std_logic := '0'; --  clk_in.clk
		clk_out_clk : out std_logic;        -- clk_out.clk
		reset_reset : in  std_logic := '0'  --   reset.reset
	);
end entity clock50to150;

architecture rtl of clock50to150 is
	component clock50to150_pll_0 is
		port (
			refclk   : in  std_logic := 'X'; -- clk
			rst      : in  std_logic := 'X'; -- reset
			outclk_0 : out std_logic;        -- clk
			locked   : out std_logic         -- export
		);
	end component clock50to150_pll_0;

begin

	pll_0 : component clock50to150_pll_0
		port map (
			refclk   => clk_in_clk,  --  refclk.clk
			rst      => reset_reset, --   reset.reset
			outclk_0 => clk_out_clk, -- outclk0.clk
			locked   => open         -- (terminated)
		);

end architecture rtl; -- of clock50to150
